-- frame_buffer.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity frame_buffer is
	port (
		alt_vip_cl_vfb_0_control_address             : in  std_logic_vector(3 downto 0)   := (others => '0'); --       alt_vip_cl_vfb_0_control.address
		alt_vip_cl_vfb_0_control_byteenable          : in  std_logic_vector(3 downto 0)   := (others => '0'); --                               .byteenable
		alt_vip_cl_vfb_0_control_write               : in  std_logic                      := '0';             --                               .write
		alt_vip_cl_vfb_0_control_writedata           : in  std_logic_vector(31 downto 0)  := (others => '0'); --                               .writedata
		alt_vip_cl_vfb_0_control_read                : in  std_logic                      := '0';             --                               .read
		alt_vip_cl_vfb_0_control_readdata            : out std_logic_vector(31 downto 0);                     --                               .readdata
		alt_vip_cl_vfb_0_control_readdatavalid       : out std_logic;                                         --                               .readdatavalid
		alt_vip_cl_vfb_0_control_waitrequest         : out std_logic;                                         --                               .waitrequest
		alt_vip_cl_vfb_0_din_data                    : in  std_logic_vector(11 downto 0)  := (others => '0'); --           alt_vip_cl_vfb_0_din.data
		alt_vip_cl_vfb_0_din_valid                   : in  std_logic                      := '0';             --                               .valid
		alt_vip_cl_vfb_0_din_startofpacket           : in  std_logic                      := '0';             --                               .startofpacket
		alt_vip_cl_vfb_0_din_endofpacket             : in  std_logic                      := '0';             --                               .endofpacket
		alt_vip_cl_vfb_0_din_ready                   : out std_logic;                                         --                               .ready
		alt_vip_cl_vfb_0_dout_data                   : out std_logic_vector(11 downto 0);                     --          alt_vip_cl_vfb_0_dout.data
		alt_vip_cl_vfb_0_dout_valid                  : out std_logic;                                         --                               .valid
		alt_vip_cl_vfb_0_dout_startofpacket          : out std_logic;                                         --                               .startofpacket
		alt_vip_cl_vfb_0_dout_endofpacket            : out std_logic;                                         --                               .endofpacket
		alt_vip_cl_vfb_0_dout_ready                  : in  std_logic                      := '0';             --                               .ready
		alt_vip_cl_vfb_0_main_clock_clk              : in  std_logic                      := '0';             --    alt_vip_cl_vfb_0_main_clock.clk
		alt_vip_cl_vfb_0_main_reset_reset            : in  std_logic                      := '0';             --    alt_vip_cl_vfb_0_main_reset.reset
		alt_vip_cl_vfb_0_mem_clock_clk               : in  std_logic                      := '0';             --     alt_vip_cl_vfb_0_mem_clock.clk
		alt_vip_cl_vfb_0_mem_master_rd_address       : out std_logic_vector(31 downto 0);                     -- alt_vip_cl_vfb_0_mem_master_rd.address
		alt_vip_cl_vfb_0_mem_master_rd_burstcount    : out std_logic_vector(5 downto 0);                      --                               .burstcount
		alt_vip_cl_vfb_0_mem_master_rd_waitrequest   : in  std_logic                      := '0';             --                               .waitrequest
		alt_vip_cl_vfb_0_mem_master_rd_read          : out std_logic;                                         --                               .read
		alt_vip_cl_vfb_0_mem_master_rd_readdata      : in  std_logic_vector(255 downto 0) := (others => '0'); --                               .readdata
		alt_vip_cl_vfb_0_mem_master_rd_readdatavalid : in  std_logic                      := '0';             --                               .readdatavalid
		alt_vip_cl_vfb_0_mem_master_wr_address       : out std_logic_vector(31 downto 0);                     -- alt_vip_cl_vfb_0_mem_master_wr.address
		alt_vip_cl_vfb_0_mem_master_wr_burstcount    : out std_logic_vector(5 downto 0);                      --                               .burstcount
		alt_vip_cl_vfb_0_mem_master_wr_waitrequest   : in  std_logic                      := '0';             --                               .waitrequest
		alt_vip_cl_vfb_0_mem_master_wr_write         : out std_logic;                                         --                               .write
		alt_vip_cl_vfb_0_mem_master_wr_writedata     : out std_logic_vector(255 downto 0);                    --                               .writedata
		alt_vip_cl_vfb_0_mem_master_wr_byteenable    : out std_logic_vector(31 downto 0);                     --                               .byteenable
		alt_vip_cl_vfb_0_mem_reset_reset             : in  std_logic                      := '0';             --     alt_vip_cl_vfb_0_mem_reset.reset
		clk_clk                                      : in  std_logic                      := '0';             --                            clk.clk
		reset_reset_n                                : in  std_logic                      := '0'              --                          reset.reset_n
	);
end entity frame_buffer;

architecture rtl of frame_buffer is
	component frame_buffer_alt_vip_cl_vfb_0 is
		generic (
			BITS_PER_SYMBOL              : integer := 8;
			NUMBER_OF_COLOR_PLANES       : integer := 2;
			COLOR_PLANES_ARE_IN_PARALLEL : integer := 1;
			PIXELS_IN_PARALLEL           : integer := 1;
			READY_LATENCY                : integer := 1;
			MAX_WIDTH                    : integer := 1920;
			MAX_HEIGHT                   : integer := 1080;
			CLOCKS_ARE_SEPARATE          : integer := 1;
			MEM_PORT_WIDTH               : integer := 256;
			MEM_BASE_ADDR                : integer := 0;
			BURST_ALIGNMENT              : integer := 1;
			WRITE_FIFO_DEPTH             : integer := 64;
			WRITE_BURST_TARGET           : integer := 32;
			READ_FIFO_DEPTH              : integer := 64;
			READ_BURST_TARGET            : integer := 32;
			WRITER_RUNTIME_CONTROL       : integer := 0;
			READER_RUNTIME_CONTROL       : integer := 0;
			IS_FRAME_WRITER              : integer := 0;
			IS_FRAME_READER              : integer := 0;
			DROP_FRAMES                  : integer := 0;
			REPEAT_FRAMES                : integer := 0;
			DROP_REPEAT_USER             : integer := 0;
			INTERLACED_SUPPORT           : integer := 0;
			CONTROLLED_DROP_REPEAT       : integer := 0;
			DROP_INVALID_FIELDS          : integer := 0;
			MULTI_FRAME_DELAY            : integer := 1;
			IS_SYNC_MASTER               : integer := 0;
			IS_SYNC_SLAVE                : integer := 0;
			LINE_BASED_BUFFERING         : integer := 0;
			PRIORITIZE_FMAX              : integer := 0;
			USER_PACKETS_MAX_STORAGE     : integer := 0;
			MAX_SYMBOLS_PER_PACKET       : integer := 10;
			NUM_BUFFERS                  : integer := 0
		);
		port (
			main_clock                  : in  std_logic                      := 'X';             -- clk
			main_reset                  : in  std_logic                      := 'X';             -- reset
			mem_clock                   : in  std_logic                      := 'X';             -- clk
			mem_reset                   : in  std_logic                      := 'X';             -- reset
			din_data                    : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- data
			din_valid                   : in  std_logic                      := 'X';             -- valid
			din_startofpacket           : in  std_logic                      := 'X';             -- startofpacket
			din_endofpacket             : in  std_logic                      := 'X';             -- endofpacket
			din_ready                   : out std_logic;                                         -- ready
			mem_master_wr_address       : out std_logic_vector(31 downto 0);                     -- address
			mem_master_wr_burstcount    : out std_logic_vector(5 downto 0);                      -- burstcount
			mem_master_wr_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			mem_master_wr_write         : out std_logic;                                         -- write
			mem_master_wr_writedata     : out std_logic_vector(255 downto 0);                    -- writedata
			mem_master_wr_byteenable    : out std_logic_vector(31 downto 0);                     -- byteenable
			dout_data                   : out std_logic_vector(11 downto 0);                     -- data
			dout_valid                  : out std_logic;                                         -- valid
			dout_startofpacket          : out std_logic;                                         -- startofpacket
			dout_endofpacket            : out std_logic;                                         -- endofpacket
			dout_ready                  : in  std_logic                      := 'X';             -- ready
			mem_master_rd_address       : out std_logic_vector(31 downto 0);                     -- address
			mem_master_rd_burstcount    : out std_logic_vector(5 downto 0);                      -- burstcount
			mem_master_rd_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			mem_master_rd_read          : out std_logic;                                         -- read
			mem_master_rd_readdata      : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mem_master_rd_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			control_address             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- address
			control_byteenable          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			control_write               : in  std_logic                      := 'X';             -- write
			control_writedata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			control_read                : in  std_logic                      := 'X';             -- read
			control_readdata            : out std_logic_vector(31 downto 0);                     -- readdata
			control_readdatavalid       : out std_logic;                                         -- readdatavalid
			control_waitrequest         : out std_logic                                          -- waitrequest
		);
	end component frame_buffer_alt_vip_cl_vfb_0;

begin

	alt_vip_cl_vfb_0 : component frame_buffer_alt_vip_cl_vfb_0
		generic map (
			BITS_PER_SYMBOL              => 4,
			NUMBER_OF_COLOR_PLANES       => 3,
			COLOR_PLANES_ARE_IN_PARALLEL => 1,
			PIXELS_IN_PARALLEL           => 1,
			READY_LATENCY                => 1,
			MAX_WIDTH                    => 160,
			MAX_HEIGHT                   => 120,
			CLOCKS_ARE_SEPARATE          => 1,
			MEM_PORT_WIDTH               => 256,
			MEM_BASE_ADDR                => 0,
			BURST_ALIGNMENT              => 1,
			WRITE_FIFO_DEPTH             => 64,
			WRITE_BURST_TARGET           => 32,
			READ_FIFO_DEPTH              => 64,
			READ_BURST_TARGET            => 32,
			WRITER_RUNTIME_CONTROL       => 1,
			READER_RUNTIME_CONTROL       => 0,
			IS_FRAME_WRITER              => 0,
			IS_FRAME_READER              => 0,
			DROP_FRAMES                  => 0,
			REPEAT_FRAMES                => 0,
			DROP_REPEAT_USER             => 0,
			INTERLACED_SUPPORT           => 0,
			CONTROLLED_DROP_REPEAT       => 0,
			DROP_INVALID_FIELDS          => 0,
			MULTI_FRAME_DELAY            => 1,
			IS_SYNC_MASTER               => 0,
			IS_SYNC_SLAVE                => 0,
			LINE_BASED_BUFFERING         => 0,
			PRIORITIZE_FMAX              => 0,
			USER_PACKETS_MAX_STORAGE     => 0,
			MAX_SYMBOLS_PER_PACKET       => 10,
			NUM_BUFFERS                  => 2
		)
		port map (
			main_clock                  => alt_vip_cl_vfb_0_main_clock_clk,              --    main_clock.clk
			main_reset                  => alt_vip_cl_vfb_0_main_reset_reset,            --    main_reset.reset
			mem_clock                   => alt_vip_cl_vfb_0_mem_clock_clk,               --     mem_clock.clk
			mem_reset                   => alt_vip_cl_vfb_0_mem_reset_reset,             --     mem_reset.reset
			din_data                    => alt_vip_cl_vfb_0_din_data,                    --           din.data
			din_valid                   => alt_vip_cl_vfb_0_din_valid,                   --              .valid
			din_startofpacket           => alt_vip_cl_vfb_0_din_startofpacket,           --              .startofpacket
			din_endofpacket             => alt_vip_cl_vfb_0_din_endofpacket,             --              .endofpacket
			din_ready                   => alt_vip_cl_vfb_0_din_ready,                   --              .ready
			mem_master_wr_address       => alt_vip_cl_vfb_0_mem_master_wr_address,       -- mem_master_wr.address
			mem_master_wr_burstcount    => alt_vip_cl_vfb_0_mem_master_wr_burstcount,    --              .burstcount
			mem_master_wr_waitrequest   => alt_vip_cl_vfb_0_mem_master_wr_waitrequest,   --              .waitrequest
			mem_master_wr_write         => alt_vip_cl_vfb_0_mem_master_wr_write,         --              .write
			mem_master_wr_writedata     => alt_vip_cl_vfb_0_mem_master_wr_writedata,     --              .writedata
			mem_master_wr_byteenable    => alt_vip_cl_vfb_0_mem_master_wr_byteenable,    --              .byteenable
			dout_data                   => alt_vip_cl_vfb_0_dout_data,                   --          dout.data
			dout_valid                  => alt_vip_cl_vfb_0_dout_valid,                  --              .valid
			dout_startofpacket          => alt_vip_cl_vfb_0_dout_startofpacket,          --              .startofpacket
			dout_endofpacket            => alt_vip_cl_vfb_0_dout_endofpacket,            --              .endofpacket
			dout_ready                  => alt_vip_cl_vfb_0_dout_ready,                  --              .ready
			mem_master_rd_address       => alt_vip_cl_vfb_0_mem_master_rd_address,       -- mem_master_rd.address
			mem_master_rd_burstcount    => alt_vip_cl_vfb_0_mem_master_rd_burstcount,    --              .burstcount
			mem_master_rd_waitrequest   => alt_vip_cl_vfb_0_mem_master_rd_waitrequest,   --              .waitrequest
			mem_master_rd_read          => alt_vip_cl_vfb_0_mem_master_rd_read,          --              .read
			mem_master_rd_readdata      => alt_vip_cl_vfb_0_mem_master_rd_readdata,      --              .readdata
			mem_master_rd_readdatavalid => alt_vip_cl_vfb_0_mem_master_rd_readdatavalid, --              .readdatavalid
			control_address             => alt_vip_cl_vfb_0_control_address,             --       control.address
			control_byteenable          => alt_vip_cl_vfb_0_control_byteenable,          --              .byteenable
			control_write               => alt_vip_cl_vfb_0_control_write,               --              .write
			control_writedata           => alt_vip_cl_vfb_0_control_writedata,           --              .writedata
			control_read                => alt_vip_cl_vfb_0_control_read,                --              .read
			control_readdata            => alt_vip_cl_vfb_0_control_readdata,            --              .readdata
			control_readdatavalid       => alt_vip_cl_vfb_0_control_readdatavalid,       --              .readdatavalid
			control_waitrequest         => alt_vip_cl_vfb_0_control_waitrequest          --              .waitrequest
		);

end architecture rtl; -- of frame_buffer
