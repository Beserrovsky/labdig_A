--! Standard library
library IEEE;
--! Standard packages
use IEEE.std_logic_1164.ALL;
-------------------------------------------------------------------------------
-- --
-- USP, PCS3335 - Laboratório Digital A --
-- --
-------------------------------------------------------------------------------
--
-- unit name: Registrador Simples (registrador)
--
--! @brief Registrador de tamanho N
--! 
--
--! @author <Felipe Beserra (felipebeserra25@usp.br)>
--! @author <Renato Ferreira (renato.ferreiraspfc@usp.br)>
--
--! @date <01\04\2024>
--
--! @version <v0.1>
--
-------------------------------------------------------------------------------
--! @todo <Criar registrador> \n
-------------------------------------------------------------------------------

entity registrador is 
port (
    --
);
end entity;

architecture registrador_arch of registrador is	
    -- constants
    -- signals
begin
    -- processes
    -- port maps
    -- combinatory logic
end architecture;
